module Ex_Mem(
    input clk,
    //数据信号输入
    input[32-1:0] ALU_ans_Ex,
    input[32-1:0] busB_Ex,
    input[]


);

endmodule